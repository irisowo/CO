//Subject:     
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      0616086
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------
module PC_instr(
	instr,
	pc,
	PC_instr_o
    );
input 	[27:0]	instr;
input	[31:0]	pc;
output	[31:0]	PC_instr_o;
	
assign PC_instr_o = {pc[31:28], instr[27:0]};
	
endmodule

                    
                    